`timescale 1ns/1ps

module frog_chip #(
	parameter N=16
)(
	input wire clk,
	input wire rst_n,
	input wire load,
	input wire test,
	
	input wire program,
	input wire seed,

	output wire out,

	output wire [N-1:0] lfsr_test,
	output wire [N-1:0] taps_test
);

	reg [N-1:0] lfsr;
	reg [N-1:0] taps;
	
	wire feedback;
	assign feedback = ^(lfsr & taps); // XOR all together with tapped flags
	
	assign out = lfsr[0]; // out is LSB
	
	// test mode parallel read out
	assign lfsr_test = lfsr;
	assign taps_test = taps;
	
	always @(posedge clk) begin
	
		if (!rst_n) begin
			lfsr <= {N{1'b0}};
            taps <= {N{1'b0}};
		end
	
		else if (load) begin
			taps <= {program, taps[N-1:1]};
			lfsr <= {seed, lfsr[N-1:1]};
		end
		
		else if (test) begin
			taps <= {N{1'b0}}; // 0 out taps
			lfsr <= {1'b0, lfsr[N-1:1]}; // shift out
		end
		
		// enable states is when we are not in load, reset, or test
		else begin
			lfsr <= {feedback, lfsr[N-1:1]};
		end
	
	end

endmodule


